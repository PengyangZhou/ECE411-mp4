/* This is the Reorder Buffer for precise exception. */