/* This is our comparator. */