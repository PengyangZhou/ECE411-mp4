/* This is the ALU of our processor. */