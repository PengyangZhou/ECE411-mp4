/* This is the testbench for CPU */

module cpu_tb ();


    
endmodule