/* This is the parametrized reservation station. */

import rv32i_types::*;

module rs #(
    parameter DATA_WIDTH = 32,
    parameter TAG_WIDTH = 4,
    parameter TAG = 0   /* the tag of this reservation station entry */
    /* and so on... */
)(
    /* ports */
);
    
endmodule