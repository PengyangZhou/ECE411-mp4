/* This is the address unit for calculating effective address */