/* This is the load buffer, containing 5 reservation stations */