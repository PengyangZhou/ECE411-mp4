/* This is decoder. */