/* This is the parametrized regfile of our processor. */